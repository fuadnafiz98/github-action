CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 390 30 90 10
176 80 1916 912
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
88
8 2-In OR~
219 2617 1077 0 1 22
0 0
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U14A
25 -7 53 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6548 0 0
2
44152.8 1
0
14 Logic Display~
6 2619 1142 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L34
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9326 0 0
2
44152.8 0
0
14 Logic Display~
6 2505 1224 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L36
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5634 0 0
2
44152.8 0
0
14 Logic Display~
6 2583 1229 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7902 0 0
2
44152.8 0
0
14 Logic Display~
6 2542 1230 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L33
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6805 0 0
2
44152.8 1
0
8 2-In OR~
219 2534 1164 0 1 22
0 0
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U8D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
6198 0 0
2
44152.8 0
0
14 Logic Display~
6 2372 1178 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L32
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9216 0 0
2
44152.8 0
0
9 Inverter~
13 2368 1051 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U13A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 13 0
1 U
9719 0 0
2
44152.8 1
0
9 2-In AND~
219 2371 973 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U12D
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3781 0 0
2
44152.8 0
0
14 Logic Display~
6 2293 1181 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L31
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8277 0 0
2
44152.8 0
0
9 Inverter~
13 2282 1052 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
3457 0 0
2
44152.8 2
0
9 2-In AND~
219 2288 976 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U12C
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
3796 0 0
2
44152.8 1
0
8 2-In OR~
219 2291 1116 0 1 22
0 0
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U8C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
6904 0 0
2
44152.8 0
0
14 Logic Display~
6 2174 1187 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L30
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8602 0 0
2
44152.8 0
0
9 2-In AND~
219 2148 982 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U12B
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3607 0 0
2
44152.8 2
0
8 2-In OR~
219 2170 1062 0 1 22
0 0
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U8B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
9456 0 0
2
44152.8 1
0
9 2-In AND~
219 2205 980 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U12A
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3348 0 0
2
44152.8 0
0
14 Logic Display~
6 2030 1204 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L29
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7418 0 0
2
44152.8 1
0
9 Inverter~
13 2027 1088 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
3281 0 0
2
44152.8 0
0
9 Inverter~
13 1951 1087 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
3613 0 0
2
44152.8 0
0
14 Logic Display~
6 1954 1203 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L28
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9506 0 0
2
44152.8 1
0
9 2-In AND~
219 1953 981 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U11D
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
6773 0 0
2
44152.8 0
0
14 Logic Display~
6 1861 1198 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L27
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8799 0 0
2
44152.8 0
0
9 2-In AND~
219 1860 982 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U11C
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7433 0 0
2
44152.8 0
0
9 2-In AND~
219 1729 984 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U11B
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6183 0 0
2
44152.8 0
0
14 Logic Display~
6 1621 1222 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L26
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5243 0 0
2
44152.8 4
0
9 Inverter~
13 1618 1158 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
3217 0 0
2
44152.8 3
0
8 3-In OR~
219 1617 1075 0 1 22
0 0
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U7C
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 7 0
1 U
998 0 0
2
44152.8 2
0
9 2-In AND~
219 1660 983 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U11A
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
9272 0 0
2
44152.8 1
0
9 2-In AND~
219 1587 982 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U9D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3327 0 0
2
44152.8 0
0
14 Logic Display~
6 1439 1225 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L25
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
466 0 0
2
44152.8 4
0
9 Inverter~
13 1436 1161 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
6854 0 0
2
44152.8 3
0
8 3-In OR~
219 1435 1078 0 1 22
0 0
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U7B
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
7745 0 0
2
44152.8 2
0
9 2-In AND~
219 1478 986 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U9C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
5764 0 0
2
44152.8 1
0
9 2-In AND~
219 1405 985 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U9B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
5379 0 0
2
44152.8 0
0
14 Logic Display~
6 1298 1159 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L24
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7186 0 0
2
44152.8 0
0
9 Inverter~
13 1295 1073 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U10A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
9136 0 0
2
44152.8 0
0
9 2-In AND~
219 1300 987 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U9A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7143 0 0
2
44152.8 0
0
14 Logic Display~
6 1166 1207 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L23
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9634 0 0
2
44152.8 0
0
9 Inverter~
13 1163 1143 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3661 0 0
2
44152.8 0
0
8 2-In OR~
219 1163 1067 0 1 22
0 0
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U8A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4323 0 0
2
44152.8 0
0
9 2-In AND~
219 1198 985 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U6D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
9804 0 0
2
44152.8 0
0
9 2-In AND~
219 1141 987 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U6C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3981 0 0
2
44152.8 0
0
14 Logic Display~
6 980 1238 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L22
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9102 0 0
2
44152.8 0
0
9 Inverter~
13 977 1174 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
6812 0 0
2
44152.8 0
0
8 3-In OR~
219 976 1080 0 1 22
0 0
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U7A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
6462 0 0
2
44152.8 0
0
9 2-In AND~
219 1019 999 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
5184 0 0
2
44152.8 0
0
9 2-In AND~
219 946 998 0 1 22
0 0
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9835 0 0
2
44152.8 0
0
14 Logic Display~
6 839 1227 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L21
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8927 0 0
2
44152.8 0
0
14 Logic Display~
6 759 1224 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L13
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3701 0 0
2
44152.8 0
0
14 Logic Display~
6 2597 878 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L20
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5444 0 0
2
44152.8 0
0
14 Logic Display~
6 2592 803 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L19
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4858 0 0
2
44152.8 0
0
14 Logic Display~
6 2592 733 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L18
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4290 0 0
2
44152.8 0
0
14 Logic Display~
6 2595 679 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L17
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4394 0 0
2
44152.8 0
0
14 Logic Display~
6 2587 604 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7544 0 0
2
44152.8 0
0
14 Logic Display~
6 2589 564 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L15
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5696 0 0
2
44152.8 0
0
14 Logic Display~
6 2590 500 0 1 2
10 0
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L14
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5601 0 0
2
44152.8 0
0
9 4-In AND~
219 693 883 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U5A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
4406 0 0
2
44152.8 0
0
9 4-In AND~
219 692 805 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U4B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 4 0
1 U
882 0 0
2
44152.8 0
0
9 4-In AND~
219 693 738 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
3359 0 0
2
44152.8 0
0
9 4-In AND~
219 691 680 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U3B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 3 0
1 U
4933 0 0
2
44152.8 0
0
9 4-In AND~
219 696 619 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
9209 0 0
2
44152.8 0
0
9 4-In AND~
219 690 564 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
7797 0 0
2
44152.8 0
0
9 4-In AND~
219 686 498 0 1 22
0 0
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
6403 0 0
2
44152.8 0
0
13 Logic Switch~
5 524 400 0 1 11
0 0
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3709 0 0
2
44152.8 3
0
14 Logic Display~
6 524 977 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L12
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9784 0 0
2
44152.8 2
0
9 Inverter~
13 550 436 0 1 22
0 0
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6816 0 0
2
44152.8 1
0
14 Logic Display~
6 577 976 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L11
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7493 0 0
2
44152.8 0
0
13 Logic Switch~
5 437 399 0 1 11
0 0
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5587 0 0
2
44152.8 3
0
14 Logic Display~
6 437 976 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L10
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5642 0 0
2
44152.8 2
0
9 Inverter~
13 463 435 0 1 22
0 0
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3577 0 0
2
44152.8 1
0
14 Logic Display~
6 490 975 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3255 0 0
2
44152.8 0
0
13 Logic Switch~
5 350 399 0 1 11
0 0
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
345 0 0
2
44152.8 3
0
14 Logic Display~
6 350 976 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3918 0 0
2
44152.8 2
0
9 Inverter~
13 376 435 0 1 22
0 0
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3469 0 0
2
44152.8 1
0
14 Logic Display~
6 403 975 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4242 0 0
2
44152.8 0
0
14 Logic Display~
6 310 976 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4467 0 0
2
44152.8 0
0
9 Inverter~
13 283 436 0 1 22
0 0
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9394 0 0
2
44152.8 0
0
14 Logic Display~
6 257 977 0 1 2
10 0
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3767 0 0
2
44152.8 3
0
13 Logic Switch~
5 257 400 0 1 11
0 0
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7988 0 0
2
44152.8 0
0
14 Logic Display~
6 2319 258 0 1 2
10 0
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3128 0 0
2
44152.8 0
0
14 Logic Display~
6 2317 220 0 1 2
10 0
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9600 0 0
2
44152.8 0
0
14 Logic Display~
6 2313 186 0 1 2
10 0
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
464 0 0
2
44152.8 0
0
14 Logic Display~
6 2311 147 0 1 2
10 0
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3575 0 0
2
44152.8 0
0
13 Logic Switch~
5 330 262 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
872 0 0
2
44152.8 0
0
13 Logic Switch~
5 327 226 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5627 0 0
2
44152.8 0
0
13 Logic Switch~
5 327 190 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
35 0 0
2
44152.8 0
0
13 Logic Switch~
5 327 157 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6481 0 0
2
44152.8 0
0
128
0 1 0 0 0 0 0 0 1 15 0 3
2371 1019
2629 1019
2629 1061
0 2 0 0 0 0 0 0 1 18 0 3
2285 1009
2611 1009
2611 1061
3 1 0 0 0 0 0 1 2 0 0 3
2620 1107
2619 1107
2619 1128
0 1 0 0 0 0 0 0 6 14 0 3
2372 1083
2546 1083
2546 1148
2 2 0 0 0 0 0 11 6 0 0 3
2285 1070
2528 1070
2528 1148
3 1 0 0 0 0 0 6 4 0 0 3
2537 1194
2583 1194
2583 1215
3 1 0 0 0 0 0 6 5 0 0 3
2537 1194
2542 1194
2542 1216
3 1 0 0 0 0 0 6 3 0 0 3
2537 1194
2505 1194
2505 1210
0 1 0 0 0 0 0 0 12 10 0 3
2378 893
2295 893
2295 954
0 1 0 0 0 0 0 0 9 126 0 4
2257 224
2257 450
2378 450
2378 951
2 0 0 0 0 0 0 9 0 0 81 2
2360 951
2360 679
2 0 0 0 0 0 0 12 0 0 81 2
2277 954
2277 679
0 1 0 0 0 0 0 0 13 15 0 3
2371 1027
2303 1027
2303 1100
2 1 0 0 0 0 0 8 7 0 0 3
2371 1069
2372 1069
2372 1164
3 1 0 0 0 0 0 9 8 0 0 3
2369 996
2371 996
2371 1033
3 1 0 0 0 0 0 13 10 0 0 3
2294 1146
2293 1146
2293 1167
2 2 0 0 0 0 0 11 13 0 0 2
2285 1070
2285 1100
3 1 0 0 0 0 0 12 11 0 0 3
2286 999
2285 999
2285 1034
0 1 0 0 0 0 0 0 15 20 0 3
2212 621
2155 621
2155 960
1 0 0 0 0 0 0 17 0 0 125 2
2212 958
2212 262
2 0 0 0 0 0 0 17 0 0 81 2
2194 958
2194 679
2 0 0 0 0 0 0 15 0 0 82 2
2137 960
2137 607
3 1 0 0 0 0 0 16 14 0 0 3
2173 1092
2174 1092
2174 1173
3 1 0 0 0 0 0 17 16 0 0 4
2203 1003
2203 1016
2182 1016
2182 1046
3 2 0 0 0 0 0 15 16 0 0 4
2146 1005
2146 1017
2164 1017
2164 1046
0 1 0 0 0 0 0 0 19 127 0 2
2030 190
2030 1070
2 1 0 0 0 0 0 19 18 0 0 2
2030 1106
2030 1190
0 1 0 0 0 0 0 0 22 35 0 3
1733 904
1960 904
1960 959
2 0 0 0 0 0 0 22 0 0 83 2
1942 959
1942 563
2 1 0 0 0 0 0 20 21 0 0 2
1954 1105
1954 1189
3 1 0 0 0 0 0 22 20 0 0 3
1951 1004
1954 1004
1954 1069
0 1 0 0 0 0 0 0 24 37 0 3
1667 898
1867 898
1867 960
2 0 0 0 0 0 0 24 0 0 79 2
1849 960
1849 805
3 1 0 0 0 0 0 24 23 0 0 4
1858 1005
1858 1178
1861 1178
1861 1184
0 1 0 0 0 0 0 0 25 39 0 3
1594 904
1736 904
1736 962
2 0 0 0 0 0 0 25 0 0 81 2
1718 962
1718 679
0 1 0 0 0 0 0 0 29 55 0 4
1306 899
1306 898
1667 898
1667 961
2 0 0 0 0 0 0 29 0 0 82 2
1649 961
1649 607
1 0 0 0 0 0 0 30 0 0 46 3
1594 960
1594 904
1485 904
2 0 0 0 0 0 0 30 0 0 84 2
1576 960
1576 498
2 1 0 0 0 0 0 27 26 0 0 2
1621 1176
1621 1208
4 1 0 0 0 0 0 28 27 0 0 4
1620 1105
1620 1132
1621 1132
1621 1140
1 3 0 0 0 0 0 28 25 0 0 4
1629 1059
1629 1020
1727 1020
1727 1007
2 3 0 0 0 0 0 28 29 0 0 4
1620 1060
1620 1014
1658 1014
1658 1006
3 3 0 0 0 0 0 28 30 0 0 4
1611 1059
1611 1013
1585 1013
1585 1005
1 0 0 0 0 0 0 34 0 0 48 3
1485 964
1485 903
1412 903
2 0 0 0 0 0 0 34 0 0 83 2
1467 964
1467 564
1 0 0 0 0 0 0 35 0 0 125 2
1412 963
1412 262
2 0 0 0 0 0 0 35 0 0 84 2
1394 963
1394 498
3 0 0 0 0 0 0 33 0 0 76 3
1429 1062
1429 1048
839 1048
2 3 0 0 0 0 0 33 35 0 0 4
1438 1063
1438 1016
1403 1016
1403 1008
1 3 0 0 0 0 0 33 34 0 0 4
1447 1062
1447 1017
1476 1017
1476 1009
2 1 0 0 0 0 0 32 31 0 0 2
1439 1179
1439 1211
4 1 0 0 0 0 0 33 32 0 0 4
1438 1108
1438 1135
1439 1135
1439 1143
0 1 0 0 0 0 0 0 38 63 0 3
1187 899
1307 899
1307 965
2 0 0 0 0 0 0 38 0 0 80 2
1289 965
1289 738
2 1 0 0 0 0 0 37 36 0 0 2
1298 1091
1298 1145
3 1 0 0 0 0 0 38 37 0 0 2
1298 1010
1298 1055
2 1 0 0 0 0 0 40 39 0 0 2
1166 1161
1166 1193
3 1 0 0 0 0 0 41 40 0 0 2
1166 1097
1166 1125
3 1 0 0 0 0 0 42 41 0 0 3
1196 1008
1175 1008
1175 1051
3 2 0 0 0 0 0 43 41 0 0 3
1139 1010
1157 1010
1157 1051
2 0 0 0 0 0 0 42 0 0 65 3
1187 963
1187 899
1148 899
0 1 0 0 0 0 0 0 42 83 0 2
1205 564
1205 963
1 0 0 0 0 0 0 43 0 0 126 2
1148 965
1148 226
2 0 0 0 0 0 0 43 0 0 84 2
1130 965
1130 498
1 2 0 0 0 0 0 44 45 0 0 2
980 1224
980 1192
1 4 0 0 0 0 0 45 46 0 0 3
980 1156
979 1156
979 1110
3 0 0 0 0 0 0 46 0 0 77 5
970 1064
970 1037
780 1037
780 1036
759 1036
3 1 0 0 0 0 0 47 46 0 0 3
1017 1022
988 1022
988 1064
3 2 0 0 0 0 0 48 46 0 0 3
944 1021
979 1021
979 1065
0 1 0 0 0 0 0 0 47 74 0 3
953 921
1026 921
1026 977
2 0 0 0 0 0 0 47 0 0 83 2
1008 977
1008 564
1 0 0 0 0 0 0 48 0 0 126 2
953 976
953 226
2 0 0 0 0 0 0 48 0 0 84 2
935 976
935 498
0 1 0 0 0 0 0 0 49 127 0 2
839 190
839 1213
0 1 0 0 0 0 0 0 50 128 0 2
759 157
759 1210
5 1 0 0 0 0 0 58 51 0 0 4
714 883
729 883
729 881
2582 881
5 1 0 0 0 0 0 59 52 0 0 4
713 805
1849 805
1849 806
2577 806
5 1 0 0 0 0 0 60 53 0 0 4
714 738
1639 738
1639 736
2577 736
5 1 0 0 0 0 0 61 54 0 0 5
712 680
1620 680
1620 679
2580 679
2580 682
5 1 0 0 0 16 0 62 55 0 0 4
717 619
727 619
727 607
2572 607
5 1 0 0 0 0 0 63 56 0 0 6
711 564
1625 564
1625 563
1942 563
1942 567
2574 567
5 1 0 0 0 0 0 64 57 0 0 4
707 498
1576 498
1576 503
2575 503
4 0 0 0 0 0 0 58 0 0 113 2
669 897
577 897
3 0 0 0 0 0 0 58 0 0 118 2
669 888
437 888
2 0 0 0 0 0 0 58 0 0 119 2
669 879
403 879
1 0 0 0 0 0 0 58 0 0 124 4
669 870
262 870
262 871
257 871
4 0 0 0 0 0 0 59 0 0 115 2
668 819
524 819
3 0 0 0 0 0 0 59 0 0 116 2
668 810
490 810
2 0 0 0 0 0 0 59 0 0 119 2
668 801
403 801
1 0 0 0 0 0 0 59 0 0 124 4
668 792
262 792
262 793
257 793
4 0 0 0 0 0 0 60 0 0 115 2
669 752
524 752
3 0 0 0 0 0 0 60 0 0 118 2
669 743
437 743
2 0 0 0 0 0 0 60 0 0 121 2
669 734
350 734
1 0 0 0 0 0 0 60 0 0 122 2
669 725
310 725
4 0 0 0 0 0 0 61 0 0 113 4
667 694
582 694
582 695
577 695
3 0 0 0 0 0 0 61 0 0 118 2
667 685
437 685
2 0 0 0 0 0 0 61 0 0 121 2
667 676
350 676
1 0 0 0 0 0 0 61 0 0 122 2
667 667
310 667
4 0 0 0 0 0 0 62 0 0 115 2
672 633
524 633
3 0 0 0 0 0 0 62 0 0 118 2
672 624
437 624
2 0 0 0 0 0 0 62 0 0 119 4
672 615
408 615
408 616
403 616
1 0 0 0 0 0 0 62 0 0 122 2
672 606
310 606
4 0 0 0 0 0 0 63 0 0 115 4
666 578
529 578
529 579
524 579
3 0 0 0 0 0 0 63 0 0 116 2
666 569
490 569
2 0 0 0 0 0 0 63 0 0 119 2
666 560
403 560
1 0 0 0 0 0 0 63 0 0 122 2
666 551
310 551
4 0 0 0 0 0 0 64 0 0 113 2
662 512
577 512
3 0 0 0 0 0 0 64 0 0 116 2
662 503
490 503
2 0 0 0 0 0 0 64 0 0 119 2
662 494
403 494
1 0 0 0 0 0 0 64 0 0 122 4
662 485
315 485
315 486
310 486
2 1 0 0 0 0 0 67 68 0 0 3
571 436
577 436
577 962
1 0 0 0 0 0 0 67 0 0 115 2
535 436
524 436
1 1 0 0 0 0 0 65 66 0 0 2
524 412
524 963
2 1 0 0 0 0 0 71 72 0 0 3
484 435
490 435
490 961
1 0 0 0 0 0 0 71 0 0 118 2
448 435
437 435
1 1 0 0 0 0 0 69 70 0 0 2
437 411
437 962
2 1 0 0 0 0 0 75 76 0 0 3
397 435
403 435
403 961
1 0 0 0 0 0 0 75 0 0 121 2
361 435
350 435
1 1 0 0 0 0 0 73 74 0 0 2
350 411
350 962
2 1 0 0 0 0 0 78 77 0 0 3
304 436
310 436
310 962
1 0 0 0 0 0 0 78 0 0 124 2
268 436
257 436
1 1 0 0 0 0 0 80 79 0 0 2
257 412
257 963
1 1 0 0 0 0 0 85 81 0 0 2
342 262
2303 262
1 1 0 0 0 0 0 86 82 0 0 4
339 226
1148 226
1148 224
2301 224
1 1 0 0 0 0 0 87 83 0 0 2
339 190
2297 190
1 1 0 0 0 0 0 88 84 0 0 4
339 157
759 157
759 151
2295 151
28
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2607 1166 2642 1190
2612 1170 2636 1186
3 CIn
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2583 1247 2610 1271
2588 1251 2604 1267
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2540 1278 2567 1302
2545 1282 2561 1298
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2499 1252 2526 1276
2504 1256 2520 1272
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2367 1203 2402 1227
2372 1207 2396 1223
3 Lo'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2285 1211 2312 1235
2290 1215 2306 1231
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2176 1196 2203 1220
2181 1200 2197 1216
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2032 1251 2067 1275
2037 1255 2061 1271
3 Li'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1949 1229 1984 1253
1954 1233 1978 1249
3 Lb'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1844 1222 1871 1246
1849 1226 1865 1242
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1617 1253 1652 1277
1622 1257 1646 1273
3 LA'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1425 1264 1460 1288
1430 1268 1454 1284
3 CE'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1295 1186 1322 1210
1300 1190 1316 1206
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1155 1237 1190 1261
1160 1241 1184 1257
3 Ei'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
978 1262 1013 1286
983 1266 1007 1282
3 LM'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
833 1246 860 1270
838 1250 854 1266
2 CP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
748 1256 775 1280
753 1260 769 1276
2 EP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
711 780 746 804
716 784 740 800
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
711 854 746 878
716 858 740 874
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
712 711 747 735
717 715 741 731
3 JMP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
714 658 749 682
719 662 743 678
3 INR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
720 588 755 612
725 592 749 608
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
710 542 745 566
715 546 739 562
3 LDB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
705 481 740 505
710 485 734 501
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
279 247 306 271
284 251 300 267
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
278 212 305 236
283 216 299 232
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
277 179 304 203
282 183 298 199
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
275 146 302 170
280 150 296 166
2 T1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
